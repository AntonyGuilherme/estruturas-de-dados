-- Code your testbench here
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY TESTES_EXERCICIO5 IS
END TESTES_EXERCICIO5;

ARCHITECTURE TESTE_COMPORTAMENTAL OF TESTES_EXERCICIO5 IS

    COMPONENT FUNCAO_X IS

        PORT (
            ENTRADA_X : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			SAIDA_FUNCAO : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
        );

    END COMPONENT FUNCAO_X;

	SIGNAL ENTRADA_X : STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL SAIDA_FUNCAO : STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
    INSTANCIA_TESTE : FUNCAO_X PORT MAP(ENTRADA_X, SAIDA_FUNCAO);
    ENTRADA_X <= "0000",
        "0110" AFTER 10 ns,
        "1111" AFTER 20 ns,
        "0000" AFTER 50 ns;

END TESTE_COMPORTAMENTAL;