-- library declaration
LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

-- entity
ENTITY FUNCAO_X IS

    PORT (
        ENTRADA_X : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
        SAIDA_FUNCAO : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
    );

END FUNCAO_X;

-- architecture
ARCHITECTURE COMPORTAMENTAL OF FUNCAO_X IS

    SIGNAL MULTIPLICACAO_X_NOT_X : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

    MULTIPLICACAO_X_NOT_X <= STD_LOGIC_VECTOR((unsigned(ENTRADA_X) * unsigned(NOT(ENTRADA_X))));
    SAIDA_FUNCAO <= STD_LOGIC_VECTOR(unsigned(MULTIPLICACAO_X_NOT_X) SLL 1);

END COMPORTAMENTAL;